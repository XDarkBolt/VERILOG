/////////////////////////////////////////
//					FREQ_DIV						//
/////////////////////////////////////////

module FREQ_DIV ( clk , clk0 );

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//SETTINGS

parameter	DIV	= 12;

//SETTINGS				
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

input clk;

output reg clk0;

/////////////////////////////////////////

reg [DIV:0] counter;

/////////////////////////////////////////

always @( posedge clk )
begin
	counter <= counter + 1;
end

/////////////////////////////////////////

always
begin
	clk0 <= counter[DIV];
end

/////////////////////////////////////////

endmodule

/////////////////////////////////////////